// DSCH 3.9
// 3/25/2025 6:17:30 PM
// E:\mos\BOOTG;S\stage1.sch

module stage1( in36,multiplicand_0,multiplier_4,acc1,in37,acc0,multiplier_7,acc2,
 multiplier_6,multiplier_5,multiplier_3,multiplier_0,acc7,multiplicand_7,multiplier_2,multiplier_1,
 multiplicand_6,multiplicand_5,acc6,multiplicand_4,multiplicand_2,acc4,acc5,multiplicand_1,
 multiplicand_3,acc3,in27,nxt0,nxt6,nxt2,nxt5,nxt3,
 nxt4,nxt1,nxt7,nxt_acc7,nxt_acc4,nxt_acc1,nxt_acc2,nxt_acc3,
 nxt_acc0,nxt_acc5,nxt_acc6);
 input in36,multiplicand_0,multiplier_4,acc1,in37,acc0,multiplier_7,acc2;
 input multiplier_6,multiplier_5,multiplier_3,multiplier_0,acc7,multiplicand_7,multiplier_2,multiplier_1;
 input multiplicand_6,multiplicand_5,acc6,multiplicand_4,multiplicand_2,acc4,acc5,multiplicand_1;
 input multiplicand_3,acc3,in27;
 output nxt0,nxt6,nxt2,nxt5,nxt3,nxt4,nxt1,nxt7;
 output nxt_acc7,nxt_acc4,nxt_acc1,nxt_acc2,nxt_acc3,nxt_acc0,nxt_acc5,nxt_acc6;
 wire w2,w4,w13,w14,w15,w16,w17,w18;
 wire w19,w20,w22,w23,w24,w25,w26,w27;
 wire w28,w29,w30,w31,w32,w33,w34,w35;
 wire w36,w37,w38,w39,w40,w41,w42,w43;
 wire w44,w45,w46,w47,w48,w49,w50,w67;
 wire w68,w69,w70,w71,w72,w73,w74,w75;
 wire w76,w77,w78,w80,w81,w82,w83,w84;
 wire w85,w86,w87,w88,w89,w90,w91,w92;
 wire w93,w94,w95,w96,w97,w106,w115,w116;
 wire w117,w118,w119,w120,w121,w122,w123,w124;
 wire w125,w126,w127,w128,w129,w130,w131,w132;
 wire w133,w134,w135,w136,w137,w138,w139,w140;
 wire w141,w142,w143,w144,w145,w146,w147,w148;
 wire w149,w150,w151,w152,w153,w154,w155,w156;
 wire w157,w158,w159,w160,w161,w162,w163,w164;
 wire w165,w166,w167,w168,w169,w170,w171,w172;
 wire w173,w174,w175,w176,w177,w178,w179,w180;
 wire w181,w182,w183,w184,w185,w186,w187,w188;
 wire w189,w190,w191,w192,w193,w194,w195,w196;
 wire w197,w198,w199,w200,w201,w202,w203,w204;
 wire w205,w206,w207,w208,w209,w210,w211,w212;
 wire w213,w214,w215,w216,w217,w218,w219,w220;
 wire w221,w222,w223,w224,w225,w226,w227,w228;
 wire w229,w230,w231,w232,w233,w234,w235,w236;
 wire w237,w238,w239,w240,w241,w242,w243,w244;
 wire w245,w246,w247,w248,w249,w250,w251,w252;
 wire w253,w254,w255,w256,w257,w258,w259,w260;
 wire w261,w262,w263,w264,w265,w266,w267,w268;
 wire w269,w270,w271,w272,w273,w274,w275,w276;
 wire w277,w278,w279,w280,w281,w282,w283,w284;
 wire w285,w286,w287,w288,w289,w290,w291,w292;
 wire w293,w294,w295,w296,w297,w298,w299,w300;
 wire w301,w302,w303,w304,w305,w306,w307,w308;
 wire w309,w310,w311,w312,w313,w314,w315,w316;
 wire w317,w318,w319,w320,w321,w322,w323,w324;
 wire w325,w326,w327,w328,w329,w330,w331,w332;
 wire w333,w334,w335,w336,w337,w338,w339,w340;
 wire w341,w342,w343,w344,w345,w346,w347,w348;
 wire w349,w350,w351,w352,w353,w354,w355,w356;
 wire w357,w358,w359,w360,w361,w362,w363,w364;
 wire w365,w366,w367,w368,w369,w370,w371,w372;
 wire w373,w374,w375,w376,w377,w378,w379,w380;
 wire w381,w382,w383,w384,w385,w386,w387,w388;
 wire w389,w390,w391,w392,w393,w394,w395,w396;
 wire w397,w398,w399,w400,w401,w402,w403,w404;
 wire w405,w406,w407,w408,w409,w410,w411,w412;
 wire w413,w414,w415,w416,w417,w418,w419,w420;
 wire w421,w422,w423,w424,w425,w426,w427,w428;
 wire w429,w430,w431,w432,w433,w434,w435,w436;
 wire w437,w438,w439,w440,w441,w442,w443,w444;
 wire w445,w446,w447,w448,w449,w450,w451,w452;
 wire w453,w454,w455,w456,w457,w458,w459,w460;
 wire w461,w462,w463,w464,w465,w466,w467,w468;
 wire w469,w470,w471,w472,w473,w474,w475,w476;
 wire w477,w478,w479,w480,w481,w482,w483,w484;
 wire w485,w486,w487,w488,w489,w490,w491,w492;
 wire w493,w494,w495,w496,w497,w498,w499,w500;
 wire w501,w502,w503,w504,w505,w506,w507,w508;
 wire w509,w510,w511,w512,w513;
 dreg #(12) dreg_1_1(w13,w117,w115,w116,w4);
 not #(8) inv_2_2(w118,w2);
 or #(8) or2_3_3(w115,w119,w120);
 and #(8) and2_4_4(w120,w118,w14);
 and #(8) and2_5_5(w119,w2,acc7);
 dreg #(12) dreg_6_6(w14,w123,w121,w122,w4);
 not #(8) inv_7_7(w124,w2);
 or #(8) or2_8_8(w121,w125,w126);
 and #(8) and2_9_9(w126,w124,w15);
 and #(8) and2_10_10(w125,w2,acc6);
 dreg #(12) dreg_11_11(w15,w129,w127,w128,w4);
 not #(8) inv_12_12(w130,w2);
 or #(8) or2_13_13(w127,w131,w132);
 and #(8) and2_14_14(w132,w130,w16);
 and #(8) and2_15_15(w131,w2,acc5);
 dreg #(12) dreg_16_16(w16,w135,w133,w134,w4);
 not #(8) inv_17_17(w136,w2);
 or #(8) or2_18_18(w133,w137,w138);
 and #(8) and2_19_19(w138,w136,w17);
 and #(8) and2_20_20(w137,w2,acc4);
 dreg #(12) dreg_21_21(w17,w141,w139,w140,w4);
 not #(8) inv_22_22(w142,w2);
 or #(8) or2_23_23(w139,w143,w144);
 and #(8) and2_24_24(w145,w2,acc0);
 and #(8) and2_25_25(w147,w146,in37);
 or #(8) or2_26_26(w148,w145,w147);
 not #(8) inv_27_27(w146,w2);
 and #(8) and2_28_28(w144,w142,w18);
 and #(8) and2_29_29(w143,w2,acc3);
 dreg #(12) dreg_30_30(w18,w151,w149,w150,w4);
 dreg #(12) dreg_31_31(w20,w153,w148,w152,w4);
 and #(8) and2_32_32(w154,w2,acc1);
 and #(8) and2_33_33(w156,w155,w20);
 or #(8) or2_34_34(w157,w154,w156);
 not #(8) inv_35_35(w155,w2);
 not #(8) inv_36_36(w158,w2);
 dreg #(12) dreg_37_37(w19,w160,w157,w159,w4);
 and #(8) and2_38_38(w161,w2,acc2);
 and #(8) and2_39_39(w162,w158,w19);
 or #(8) or2_40_40(w149,w161,w162);
 dreg #(12) dreg_1_41(w32,w165,w163,w164,w24);
 not #(8) inv_2_42(w166,w22);
 or #(8) or2_3_43(w163,w167,w168);
 and #(8) and2_4_44(w168,w166,w33);
 and #(8) and2_5_45(w167,w22,w23);
 dreg #(12) dreg_6_46(w33,w171,w169,w170,w24);
 not #(8) inv_7_47(w172,w22);
 or #(8) or2_8_48(w169,w173,w174);
 and #(8) and2_9_49(w174,w172,w34);
 and #(8) and2_10_50(w173,w22,w25);
 dreg #(12) dreg_11_51(w34,w177,w175,w176,w24);
 not #(8) inv_12_52(w178,w22);
 or #(8) or2_13_53(w175,w179,w180);
 and #(8) and2_14_54(w180,w178,w35);
 and #(8) and2_15_55(w179,w22,w27);
 dreg #(12) dreg_16_56(w35,w183,w181,w182,w24);
 not #(8) inv_17_57(w184,w22);
 or #(8) or2_18_58(w181,w185,w186);
 and #(8) and2_19_59(w186,w184,w36);
 and #(8) and2_20_60(w185,w22,w26);
 dreg #(12) dreg_21_61(w36,w189,w187,w188,w24);
 not #(8) inv_22_62(w190,w22);
 or #(8) or2_23_63(w187,w191,w192);
 and #(8) and2_24_64(w193,w22,w29);
 and #(8) and2_25_65(w195,w194,in36);
 or #(8) or2_26_66(w196,w193,w195);
 not #(8) inv_27_67(w194,w22);
 and #(8) and2_28_68(w192,w190,w37);
 and #(8) and2_29_69(w191,w22,w28);
 dreg #(12) dreg_30_70(w37,w199,w197,w198,w24);
 dreg #(12) dreg_31_71(w39,w201,w196,w200,w24);
 and #(8) and2_32_72(w202,w22,w30);
 and #(8) and2_33_73(w204,w203,w39);
 or #(8) or2_34_74(w205,w202,w204);
 not #(8) inv_35_75(w203,w22);
 not #(8) inv_36_76(w206,w22);
 dreg #(12) dreg_37_77(w38,w208,w205,w207,w24);
 and #(8) and2_38_78(w209,w22,w31);
 and #(8) and2_39_79(w210,w206,w38);
 or #(8) or2_40_80(w197,w209,w210);
 not #(10) inv_1_81(w212,w211);
 nand #(21) nand2_2_82(w214,w213,w212);
 nand #(21) nand2_3_83(w215,w214,w214);
 nand #(21) nand2_4_84(w217,w211,w216);
 nand #(21) nand2_5_85(w218,w217,w217);
 nand #(27) nand2_6_86(w28,w219,w220);
 nand #(13) nand2_7_87(w219,w215,w215);
 nand #(13) nand2_8_88(w220,w218,w218);
 not #(10) inv_9_89(w216,w213);
 nand #(13) nand2_10_90(w222,w221,w221);
 nand #(13) nand2_11_91(w224,w223,w223);
 nand #(21) nand2_12_92(w223,w225,w225);
 nand #(21) nand2_13_93(w225,w226,acc3);
 nand #(21) nand2_14_94(w211,w224,w222);
 nand #(21) nand2_15_95(w221,w227,w227);
 nand #(21) nand2_16_96(w227,w40,w228);
 not #(10) inv_17_97(w228,acc3);
 not #(10) inv_18_98(w226,w40);
 nand #(21) nand2_19_99(w229,w40,acc3);
 nand #(21) nand2_20_100(w230,w229,w229);
 nand #(21) nand2_21_101(w231,w40,w213);
 nand #(21) nand2_22_102(w232,w231,w231);
 nand #(21) nand2_23_103(w233,w213,acc3);
 nand #(21) nand2_24_104(w234,w233,w233);
 nand #(13) nand2_25_105(w235,w230,w230);
 nand #(13) nand2_26_106(w236,w232,w232);
 nand #(21) nand2_27_107(w237,w236,w235);
 nand #(13) nand2_28_108(w238,w237,w237);
 nand #(13) nand2_29_109(w239,w234,w234);
 nand #(34) nand2_30_110(w45,w239,w238);
 not #(10) inv_31_111(w241,w240);
 nand #(21) nand2_32_112(w243,w242,w241);
 nand #(21) nand2_33_113(w244,w243,w243);
 nand #(21) nand2_34_114(w246,w240,w245);
 nand #(21) nand2_35_115(w247,w246,w246);
 nand #(27) nand2_36_116(w31,w248,w249);
 nand #(13) nand2_37_117(w248,w244,w244);
 nand #(13) nand2_38_118(w249,w247,w247);
 not #(10) inv_39_119(w245,w242);
 nand #(13) nand2_40_120(w251,w250,w250);
 nand #(13) nand2_41_121(w253,w252,w252);
 nand #(21) nand2_42_122(w252,w254,w254);
 nand #(21) nand2_43_123(w254,w255,acc2);
 nand #(21) nand2_44_124(w240,w253,w251);
 nand #(21) nand2_45_125(w250,w256,w256);
 nand #(21) nand2_46_126(w256,w41,w257);
 not #(10) inv_47_127(w257,acc2);
 not #(10) inv_48_128(w255,w41);
 nand #(21) nand2_49_129(w258,w41,acc2);
 nand #(21) nand2_50_130(w259,w258,w258);
 nand #(21) nand2_51_131(w260,w41,w242);
 nand #(21) nand2_52_132(w261,w260,w260);
 nand #(21) nand2_53_133(w264,w262,w263);
 nand #(21) nand2_54_134(w265,w242,acc2);
 nand #(21) nand2_55_135(w266,w265,w265);
 nand #(13) nand2_56_136(w267,w259,w259);
 nand #(13) nand2_57_137(w268,w261,w261);
 nand #(21) nand2_58_138(w269,w268,w267);
 nand #(13) nand2_59_139(w270,w269,w269);
 nand #(13) nand2_60_140(w271,w266,w266);
 nand #(35) nand2_61_141(w213,w271,w270);
 nand #(21) nand2_62_142(w272,w264,w264);
 not #(10) inv_63_143(w274,w273);
 nand #(21) nand2_64_144(w276,w275,w274);
 nand #(21) nand2_65_145(w277,w276,w276);
 nand #(21) nand2_66_146(w279,w273,w278);
 nand #(21) nand2_67_147(w280,w279,w279);
 nand #(27) nand2_68_148(w30,w281,w282);
 nand #(13) nand2_69_149(w281,w277,w277);
 nand #(13) nand2_70_150(w282,w280,w280);
 not #(10) inv_71_151(w278,w275);
 nand #(13) nand2_72_152(w284,w283,w283);
 nand #(13) nand2_73_153(w286,w285,w285);
 nand #(21) nand2_74_154(w285,w287,w287);
 nand #(21) nand2_75_155(w287,w288,acc1);
 nand #(21) nand2_76_156(w273,w286,w284);
 nand #(21) nand2_77_157(w290,w43,w289);
 nand #(21) nand2_78_158(w283,w291,w291);
 nand #(21) nand2_79_159(w291,w42,w292);
 not #(10) inv_80_160(w292,acc1);
 not #(10) inv_81_161(w288,w42);
 nand #(21) nand2_82_162(w293,w42,acc1);
 nand #(21) nand2_83_163(w294,w293,w293);
 nand #(21) nand2_84_164(w295,w42,w275);
 nand #(21) nand2_85_165(w296,w295,w295);
 nand #(21) nand2_86_166(w297,w275,acc1);
 nand #(21) nand2_87_167(w298,w297,w297);
 nand #(13) nand2_88_168(w299,w294,w294);
 nand #(13) nand2_89_169(w300,w296,w296);
 nand #(21) nand2_90_170(w301,w300,w299);
 nand #(13) nand2_91_171(w302,w301,w301);
 nand #(13) nand2_92_172(w303,w298,w298);
 nand #(35) nand2_93_173(w242,w303,w302);
 nand #(21) nand2_94_174(w304,w290,w290);
 not #(10) inv_95_175(w289,w262);
 nand #(27) nand2_96_176(w29,w305,w306);
 nand #(35) nand2_97_177(w275,w307,w308);
 nand #(13) nand2_98_178(w307,w309,w309);
 nand #(13) nand2_99_179(w308,w310,w310);
 nand #(21) nand2_100_180(w310,w311,w312);
 nand #(13) nand2_101_181(w311,w313,w313);
 nand #(13) nand2_102_182(w312,w314,w314);
 nand #(21) nand2_103_183(w309,w315,w315);
 nand #(21) nand2_104_184(w315,w43,acc0);
 nand #(21) nand2_105_185(w313,w316,w316);
 nand #(21) nand2_106_186(w316,w44,w43);
 nand #(21) nand2_107_187(w314,w317,w317);
 nand #(21) nand2_108_188(w317,w44,acc0);
 not #(10) inv_109_189(w318,w44);
 not #(10) inv_110_190(w319,acc0);
 nand #(21) nand2_111_191(w320,w44,w319);
 nand #(21) nand2_112_192(w321,w320,w320);
 nand #(21) nand2_113_193(w262,w322,w323);
 nand #(21) nand2_114_194(w324,w318,acc0);
 nand #(21) nand2_115_195(w325,w324,w324);
 nand #(13) nand2_116_196(w322,w325,w325);
 nand #(13) nand2_117_197(w323,w321,w321);
 not #(10) inv_118_198(w263,w43);
 nand #(13) nand2_119_199(w306,w272,w272);
 nand #(13) nand2_120_200(w305,w304,w304);
 not #(10) inv_1_201(w327,w326);
 nand #(21) nand2_2_202(w329,w328,w327);
 nand #(21) nand2_3_203(w330,w329,w329);
 nand #(21) nand2_4_204(w332,w326,w331);
 nand #(21) nand2_5_205(w333,w332,w332);
 nand #(27) nand2_6_206(w23,w334,w335);
 nand #(13) nand2_7_207(w334,w330,w330);
 nand #(13) nand2_8_208(w335,w333,w333);
 not #(10) inv_9_209(w331,w328);
 nand #(13) nand2_10_210(w337,w336,w336);
 nand #(13) nand2_11_211(w339,w338,w338);
 nand #(21) nand2_12_212(w338,w340,w340);
 nand #(21) nand2_13_213(w340,w341,acc7);
 nand #(21) nand2_14_214(w326,w339,w337);
 nand #(21) nand2_15_215(w336,w342,w342);
 nand #(21) nand2_16_216(w342,w46,w343);
 not #(10) inv_17_217(w343,acc7);
 not #(10) inv_18_218(w341,w46);
 nand #(21) nand2_19_219(w344,w46,acc7);
 nand #(21) nand2_20_220(w345,w344,w344);
 nand #(21) nand2_21_221(w346,w46,w328);
 nand #(21) nand2_22_222(w347,w346,w346);
 nand #(21) nand2_23_223(w348,w328,acc7);
 nand #(21) nand2_24_224(w349,w348,w348);
 nand #(13) nand2_25_225(w350,w345,w345);
 nand #(13) nand2_26_226(w351,w347,w347);
 nand #(21) nand2_27_227(w352,w351,w350);
 nand #(13) nand2_28_228(w353,w352,w352);
 nand #(13) nand2_29_229(w354,w349,w349);
 nand #(6) nand2_30_230(w50,w354,w353);
 not #(10) inv_31_231(w356,w355);
 nand #(21) nand2_32_232(w358,w357,w356);
 nand #(21) nand2_33_233(w359,w358,w358);
 nand #(21) nand2_34_234(w361,w355,w360);
 nand #(21) nand2_35_235(w362,w361,w361);
 nand #(27) nand2_36_236(w25,w363,w364);
 nand #(13) nand2_37_237(w363,w359,w359);
 nand #(13) nand2_38_238(w364,w362,w362);
 not #(10) inv_39_239(w360,w357);
 nand #(13) nand2_40_240(w366,w365,w365);
 nand #(13) nand2_41_241(w368,w367,w367);
 nand #(21) nand2_42_242(w367,w369,w369);
 nand #(21) nand2_43_243(w369,w370,acc6);
 nand #(21) nand2_44_244(w355,w368,w366);
 nand #(21) nand2_45_245(w365,w371,w371);
 nand #(21) nand2_46_246(w371,w47,w372);
 not #(10) inv_47_247(w372,acc6);
 not #(10) inv_48_248(w370,w47);
 nand #(21) nand2_49_249(w373,w47,acc6);
 nand #(21) nand2_50_250(w374,w373,w373);
 nand #(21) nand2_51_251(w375,w47,w357);
 nand #(21) nand2_52_252(w376,w375,w375);
 nand #(21) nand2_53_253(w379,w377,w378);
 nand #(21) nand2_54_254(w380,w357,acc6);
 nand #(21) nand2_55_255(w381,w380,w380);
 nand #(13) nand2_56_256(w382,w374,w374);
 nand #(13) nand2_57_257(w383,w376,w376);
 nand #(21) nand2_58_258(w384,w383,w382);
 nand #(13) nand2_59_259(w385,w384,w384);
 nand #(13) nand2_60_260(w386,w381,w381);
 nand #(35) nand2_61_261(w328,w386,w385);
 nand #(21) nand2_62_262(w387,w379,w379);
 not #(10) inv_63_263(w389,w388);
 nand #(21) nand2_64_264(w391,w390,w389);
 nand #(21) nand2_65_265(w392,w391,w391);
 nand #(21) nand2_66_266(w394,w388,w393);
 nand #(21) nand2_67_267(w395,w394,w394);
 nand #(27) nand2_68_268(w27,w396,w397);
 nand #(13) nand2_69_269(w396,w392,w392);
 nand #(13) nand2_70_270(w397,w395,w395);
 not #(10) inv_71_271(w393,w390);
 nand #(13) nand2_72_272(w399,w398,w398);
 nand #(13) nand2_73_273(w401,w400,w400);
 nand #(21) nand2_74_274(w400,w402,w402);
 nand #(21) nand2_75_275(w402,w403,acc5);
 nand #(21) nand2_76_276(w388,w401,w399);
 nand #(21) nand2_77_277(w405,w45,w404);
 nand #(21) nand2_78_278(w398,w406,w406);
 nand #(21) nand2_79_279(w406,w48,w407);
 not #(10) inv_80_280(w407,acc5);
 not #(10) inv_81_281(w403,w48);
 nand #(21) nand2_82_282(w408,w48,acc5);
 nand #(21) nand2_83_283(w409,w408,w408);
 nand #(21) nand2_84_284(w410,w48,w390);
 nand #(21) nand2_85_285(w411,w410,w410);
 nand #(21) nand2_86_286(w412,w390,acc5);
 nand #(21) nand2_87_287(w413,w412,w412);
 nand #(13) nand2_88_288(w414,w409,w409);
 nand #(13) nand2_89_289(w415,w411,w411);
 nand #(21) nand2_90_290(w416,w415,w414);
 nand #(13) nand2_91_291(w417,w416,w416);
 nand #(13) nand2_92_292(w418,w413,w413);
 nand #(35) nand2_93_293(w357,w418,w417);
 nand #(21) nand2_94_294(w419,w405,w405);
 not #(10) inv_95_295(w404,w377);
 nand #(27) nand2_96_296(w26,w420,w421);
 nand #(35) nand2_97_297(w390,w422,w423);
 nand #(13) nand2_98_298(w422,w424,w424);
 nand #(13) nand2_99_299(w423,w425,w425);
 nand #(21) nand2_100_300(w425,w426,w427);
 nand #(13) nand2_101_301(w426,w428,w428);
 nand #(13) nand2_102_302(w427,w429,w429);
 nand #(21) nand2_103_303(w424,w430,w430);
 nand #(21) nand2_104_304(w430,w45,acc4);
 nand #(21) nand2_105_305(w428,w431,w431);
 nand #(21) nand2_106_306(w431,w49,w45);
 nand #(21) nand2_107_307(w429,w432,w432);
 nand #(21) nand2_108_308(w432,w49,acc4);
 not #(10) inv_109_309(w433,w49);
 not #(10) inv_110_310(w434,acc4);
 nand #(21) nand2_111_311(w435,w49,w434);
 nand #(21) nand2_112_312(w436,w435,w435);
 nand #(21) nand2_113_313(w377,w437,w438);
 nand #(21) nand2_114_314(w439,w433,acc4);
 nand #(21) nand2_115_315(w440,w439,w439);
 nand #(13) nand2_116_316(w437,w440,w440);
 nand #(13) nand2_117_317(w438,w436,w436);
 not #(10) inv_118_318(w378,w45);
 nand #(13) nand2_119_319(w421,w387,w387);
 nand #(13) nand2_120_320(w420,w419,w419);
 xor #(29) xor2_1_321(w44,multiplicand_0,multiplier_0);
 xor #(29) xor2_2_322(w42,multiplicand_1,multiplier_1);
 xor #(29) xor2_3_323(w41,multiplicand_2,multiplier_2);
 xor #(29) xor2_4_324(w40,multiplicand_3,multiplier_3);
 xor #(29) xor2_5_325(w49,multiplicand_4,multiplier_4);
 xor #(29) xor2_6_326(w48,multiplicand_5,multiplier_5);
 xor #(29) xor2_7_327(w47,multiplicand_6,multiplier_6);
 xor #(29) xor2_8_328(w46,multiplicand_7,multiplier_7);
 dreg #(12) dreg_1_329(w70,w443,w441,w442,w68);
 not #(8) inv_2_330(w444,w67);
 or #(8) or2_3_331(w441,w445,w446);
 and #(8) and2_4_332(w446,w444,w71);
 and #(8) and2_5_333(w445,w67,acc7);
 dreg #(12) dreg_6_334(w71,w449,w447,w448,w68);
 not #(8) inv_7_335(w450,w67);
 or #(8) or2_8_336(w447,w451,w452);
 and #(8) and2_9_337(w452,w450,w72);
 and #(8) and2_10_338(w451,w67,acc6);
 dreg #(12) dreg_11_339(w72,w455,w453,w454,w68);
 not #(8) inv_12_340(w456,w67);
 or #(8) or2_13_341(w453,w457,w458);
 and #(8) and2_14_342(w458,w456,w73);
 and #(8) and2_15_343(w457,w67,acc5);
 dreg #(12) dreg_16_344(w73,w461,w459,w460,w68);
 not #(8) inv_17_345(w462,w67);
 or #(8) or2_18_346(w459,w463,w464);
 and #(8) and2_19_347(w464,w462,w74);
 and #(8) and2_20_348(w463,w67,acc4);
 dreg #(12) dreg_21_349(w74,w467,w465,w466,w68);
 not #(8) inv_22_350(w468,w67);
 or #(8) or2_23_351(w465,w469,w470);
 and #(8) and2_24_352(w471,w67,acc0);
 and #(8) and2_25_353(w473,w472,w69);
 or #(8) or2_26_354(w474,w471,w473);
 not #(8) inv_27_355(w472,w67);
 and #(8) and2_28_356(w470,w468,w75);
 and #(8) and2_29_357(w469,w67,acc3);
 dreg #(12) dreg_30_358(w75,w477,w475,w476,w68);
 dreg #(12) dreg_31_359(w77,w479,w474,w478,w68);
 and #(8) and2_32_360(w480,w67,acc1);
 and #(8) and2_33_361(w482,w481,w77);
 or #(8) or2_34_362(w483,w480,w482);
 not #(8) inv_35_363(w481,w67);
 not #(8) inv_36_364(w484,w67);
 dreg #(12) dreg_37_365(w76,w486,w483,w485,w68);
 and #(8) and2_38_366(w487,w67,acc2);
 and #(8) and2_39_367(w488,w484,w76);
 or #(8) or2_40_368(w475,w487,w488);
 nand #(13) nand2_1_369(w490,w489,acc0);
 nand #(13) nand2_2_370(w491,multiplicand_0,w489);
 nand #(21) nand2_3_371(w489,multiplicand_0,acc0);
 nand #(13) nand2_4_372(w492,w491,w490);
 not #(10) inv_5_373(w493,w492);
 and #(16) and2_6_374(w496,w494,w495);
 and #(135) and2_7_375(w78,w496,w497);
 and #(16) and2_8_376(w497,w498,w499);
 and #(16) and2_9_377(w494,w500,w501);
 and #(16) and2_10_378(w495,w502,w503);
 and #(16) and2_11_379(w498,w504,w505);
 and #(16) and2_12_380(w499,w506,w493);
 nand #(13) nand2_13_381(w508,w507,acc1);
 nand #(13) nand2_14_382(w509,multiplicand_1,w507);
 nand #(21) nand2_15_383(w507,multiplicand_1,acc1);
 nand #(13) nand2_16_384(w510,w509,w508);
 not #(10) inv_17_385(w506,w510);
 nand #(13) nand2_18_386(w512,w511,acc2);
 nand #(13) nand2_19_387(w513,multiplicand_2,w511);
 nand #(21) nand2_20_388(w511,multiplicand_2,acc2);
 nand #(13) nand2_21_389(w514,w513,w512);
 not #(10) inv_22_390(w505,w514);
 nand #(13) nand2_23_391(w516,w515,acc3);
 nand #(13) nand2_24_392(w517,multiplicand_3,w515);
 nand #(21) nand2_25_393(w515,multiplicand_3,acc3);
 nand #(13) nand2_26_394(w518,w517,w516);
 not #(10) inv_27_395(w504,w518);
 nand #(13) nand2_28_396(w520,w519,acc4);
 nand #(13) nand2_29_397(w521,multiplicand_4,w519);
 nand #(21) nand2_30_398(w519,multiplicand_4,acc4);
 nand #(13) nand2_31_399(w522,w521,w520);
 not #(10) inv_32_400(w503,w522);
 nand #(13) nand2_33_401(w524,w523,acc5);
 nand #(13) nand2_34_402(w525,multiplicand_5,w523);
 nand #(21) nand2_35_403(w523,multiplicand_5,acc5);
 nand #(13) nand2_36_404(w526,w525,w524);
 not #(10) inv_37_405(w502,w526);
 nand #(13) nand2_38_406(w528,w527,acc6);
 nand #(13) nand2_39_407(w529,multiplicand_6,w527);
 nand #(21) nand2_40_408(w527,multiplicand_6,acc6);
 nand #(13) nand2_41_409(w530,w529,w528);
 not #(10) inv_42_410(w501,w530);
 nand #(13) nand2_43_411(w532,w531,acc7);
 nand #(13) nand2_44_412(w533,multiplicand_7,w531);
 nand #(21) nand2_45_413(w531,multiplicand_7,acc7);
 nand #(13) nand2_46_414(w534,w533,w532);
 not #(10) inv_47_415(w500,w534);
 not #(10) inv_1_416(w535,w23);
 or #(16) or2_2_417(w80,w536,w537);
 and #(16) and2_3_418(w537,w32,w23);
 and #(16) and2_4_419(w536,in27,w535);
 not #(10) inv_1_420(w538,w25);
 or #(16) or2_2_421(w81,w539,w540);
 and #(16) and2_3_422(w540,w33,w25);
 and #(16) and2_4_423(w539,in27,w538);
 not #(10) inv_1_424(w541,w27);
 or #(16) or2_2_425(w82,w542,w543);
 and #(16) and2_3_426(w543,w34,w27);
 and #(16) and2_4_427(w542,in27,w541);
 not #(10) inv_1_428(w544,w26);
 or #(16) or2_2_429(w83,w545,w546);
 and #(16) and2_3_430(w546,w35,w26);
 and #(16) and2_4_431(w545,in27,w544);
 not #(10) inv_1_432(w547,w28);
 or #(16) or2_2_433(w84,w548,w549);
 and #(16) and2_3_434(w549,w36,w28);
 and #(16) and2_4_435(w548,in27,w547);
 not #(10) inv_1_436(w550,w31);
 or #(16) or2_2_437(w85,w551,w552);
 and #(16) and2_3_438(w552,w37,w31);
 and #(16) and2_4_439(w551,in27,w550);
 not #(10) inv_1_440(w553,w30);
 or #(16) or2_2_441(w86,w554,w555);
 and #(16) and2_3_442(w555,w38,w30);
 and #(16) and2_4_443(w554,in27,w553);
 not #(10) inv_1_444(w556,w29);
 or #(16) or2_2_445(w87,w557,w558);
 and #(16) and2_3_446(w558,w39,w29);
 and #(16) and2_4_447(w557,in27,w556);
 not #(10) inv_1_448(w559,acc7);
 or #(16) or2_2_449(w88,w560,w561);
 and #(16) and2_3_450(w561,w13,acc7);
 and #(16) and2_4_451(w560,in27,w559);
 not #(10) inv_1_452(w562,acc6);
 or #(16) or2_2_453(w90,w563,w564);
 and #(16) and2_3_454(w564,w14,acc6);
 and #(16) and2_4_455(w563,w89,w562);
 not #(10) inv_1_456(w565,acc5);
 or #(16) or2_2_457(w91,w566,w567);
 and #(16) and2_3_458(w567,w15,acc5);
 and #(16) and2_4_459(w566,in27,w565);
 not #(10) inv_1_460(w568,acc4);
 or #(16) or2_2_461(w92,w569,w570);
 and #(16) and2_3_462(w570,w16,acc4);
 and #(16) and2_4_463(w569,in27,w568);
 not #(10) inv_1_464(w571,acc3);
 or #(16) or2_2_465(w94,w572,w573);
 and #(16) and2_3_466(w573,w17,acc3);
 and #(16) and2_4_467(w572,w93,w571);
 not #(10) inv_1_468(w574,acc2);
 or #(16) or2_2_469(w95,w575,w576);
 and #(16) and2_3_470(w576,w18,acc2);
 and #(16) and2_4_471(w575,in27,w574);
 not #(10) inv_1_472(w577,acc1);
 or #(16) or2_2_473(w96,w578,w579);
 and #(16) and2_3_474(w579,w19,acc1);
 and #(16) and2_4_475(w578,in27,w577);
 not #(10) inv_1_476(w580,acc0);
 or #(16) or2_2_477(w97,w581,w582);
 and #(16) and2_3_478(w582,w20,acc0);
 and #(16) and2_4_479(w581,in27,w580);
 or #(15) or2_1_480(nxt7,w583,w584);
 and #(15) and2_2_481(w584,w80,w78);
 and #(15) and2_3_482(w583,w88,w585);
 and #(15) and2_4_483(w586,w97,w585);
 and #(15) and2_5_484(w587,w87,w78);
 or #(15) or2_6_485(nxt0,w586,w587);
 not #(86) inv_7_486(w585,w78);
 or #(15) or2_8_487(nxt6,w588,w589);
 and #(15) and2_9_488(w589,w81,w78);
 and #(15) and2_10_489(w588,w90,w585);
 and #(15) and2_11_490(w590,w96,w585);
 and #(15) and2_12_491(w591,w86,w78);
 or #(15) or2_13_492(nxt1,w590,w591);
 and #(15) and2_14_493(w592,w95,w585);
 and #(15) and2_15_494(w593,w85,w78);
 or #(15) or2_16_495(nxt2,w592,w593);
 and #(15) and2_17_496(w594,w94,w585);
 and #(15) and2_18_497(w595,w84,w78);
 or #(15) or2_19_498(nxt3,w594,w595);
 and #(15) and2_20_499(w596,w92,w585);
 and #(15) and2_21_500(w597,w83,w78);
 or #(15) or2_22_501(nxt4,w596,w597);
 and #(15) and2_23_502(w598,w91,w585);
 and #(15) and2_24_503(w599,w82,w78);
 or #(15) or2_25_504(nxt5,w598,w599);
 or #(15) or2_1_505(nxt_acc7,w600,w601);
 and #(15) and2_2_506(w601,w70,w78);
 and #(15) and2_3_507(w600,in27,w602);
 and #(15) and2_4_508(w603,in27,w602);
 and #(15) and2_5_509(w604,w77,w78);
 or #(15) or2_6_510(nxt_acc0,w603,w604);
 not #(86) inv_7_511(w602,w78);
 or #(15) or2_8_512(nxt_acc6,w605,w606);
 and #(15) and2_9_513(w606,w71,w78);
 and #(15) and2_10_514(w605,in27,w602);
 and #(15) and2_11_515(w607,in27,w602);
 and #(15) and2_12_516(w608,w106,w78);
 or #(15) or2_13_517(nxt_acc1,w607,w608);
 and #(15) and2_14_518(w609,in27,w602);
 and #(15) and2_15_519(w610,w75,w78);
 or #(15) or2_16_520(nxt_acc2,w609,w610);
 and #(15) and2_17_521(w611,in27,w602);
 and #(15) and2_18_522(w612,w74,w78);
 or #(15) or2_19_523(nxt_acc3,w611,w612);
 and #(15) and2_20_524(w613,in27,w602);
 and #(15) and2_21_525(w614,w73,w78);
 or #(15) or2_22_526(nxt_acc4,w613,w614);
 and #(15) and2_23_527(w615,in27,w602);
 and #(15) and2_24_528(w616,w72,w78);
 or #(15) or2_25_529(nxt_acc5,w615,w616);
endmodule

// Simulation parameters in Verilog Format
always
#100 in36=~in36;
#200 multiplicand-0=~multiplicand-0;
#400 multiplier-4=~multiplier-4;
#800 acc1=~acc1;
#1600 in37=~in37;
#3200 acc0=~acc0;
#6400 multiplier-7=~multiplier-7;
#12800 acc2=~acc2;
#25600 multiplier-6=~multiplier-6;
#51200 multiplier-5=~multiplier-5;
#51200 multiplier-3=~multiplier-3;
#51200 multiplier-0=~multiplier-0;
#51200 acc7=~acc7;
#51200 multiplicand-7=~multiplicand-7;
#51200 multiplier-2=~multiplier-2;
#51200 multiplier-1=~multiplier-1;
#51200 multiplicand-6=~multiplicand-6;
#51200 multiplicand-5=~multiplicand-5;
#51200 acc6=~acc6;
#51200 multiplicand-4=~multiplicand-4;
#51200 multiplicand-2=~multiplicand-2;
#51200 acc4=~acc4;
#51200 acc5=~acc5;
#51200 multiplicand-1=~multiplicand-1;
#51200 multiplicand-3=~multiplicand-3;
#51200 acc3=~acc3;
#51200 in27=~in27;

// Simulation parameters
// in36 CLK 1 1
// multiplicand-0 CLK 2 2
// multiplier-4 CLK 4 4
// acc1 CLK 8 8
// in37 CLK 16 16
// acc0 CLK 32 32
// multiplier-7 CLK 64 64
// acc2 CLK 128 128
// multiplier-6 CLK 256 256
// multiplier-5 CLK 512 512
// multiplier-3 CLK 1024 1024
// multiplier-0 CLK 2048 2048
// acc7 CLK 4096 4096
// multiplicand-7 CLK 8192 8192
// multiplier-2 CLK 16384 16384
// multiplier-1 CLK 32768 32768
// multiplicand-6 CLK 32768 32768
// multiplicand-5 CLK 32768 32768
// acc6 CLK 32768 32768
// multiplicand-4 CLK 32768 32768
// multiplicand-2 CLK 32768 32768
// acc4 CLK 32768 32768
// acc5 CLK 32768 32768
// multiplicand-1 CLK 32768 32768
// multiplicand-3 CLK 32768 32768
// acc3 CLK 32768 32768
// in27 CLK 32768 32768
